module top_module (input a, input b, input c, output out);//

    nand inst1 ( out, a, b, c );

endmodule
